package driver_pkg;
    import generator_pkg :: convdata;
endpackage: driver_pkg